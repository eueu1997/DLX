package CONSTANTS is
   constant STEP : integer := 4;
   constant WORD : integer := 32;
end CONSTANTS;

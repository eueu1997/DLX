package CONSTANTS is
   constant bit_data : integer := 32;
   constant bit_add : integer := 5;
end CONSTANTS;

library ieee;
use ieee.std_logic_1164.all;

entity prova_tb is
 end prova_tb;

architecture tb of prova_tbis

generic ( nbit : integer );

endcomponent;

